`timescale 1ns / 1ps

module Div(

input [3:0]x,y,
output [3:0]z

    );

assign z=x/y;



endmodule
