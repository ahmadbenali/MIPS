// Verilog test fixture created from schematic C:\AMD\first\TT.sch - Thu Oct 05 02:55:05 2023

`timescale 1ns / 1ps

module TT_TT_sch_tb();

// Inputs

// Output

// Bidirs

// Instantiate the UUT
   TT UUT (
		
   );
// Initialize Inputs
   `ifdef auto_init
       initial begin
   `endif
endmodule
