`timescale 1ns / 1ps

module HS_SL(x,y,s,B);

input x,y;
output s,B;

wire z;

xor


endmodule
