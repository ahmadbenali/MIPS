`timescale 1ns / 1ps

module FSS();


endmodule
