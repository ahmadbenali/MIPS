`timescale 1ns / 1ps

module Load_instruction(


   
);


endmodule
