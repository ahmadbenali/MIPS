`timescale 1ns / 1ps

module ShiftRightReg
#(parameter N=4)
(

input [3:0]in ,
input CLK ,
output reg [3:0]Q
    );





endmodule
